module or2(a, b, y);
    input a, b;     // entradas
    output y;       // saida

    or(y, a, b);    // porta logica OR
    
endmodule