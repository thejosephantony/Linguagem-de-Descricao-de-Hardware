module inv(a, y);  // inversor
    input a;        // entrada
    output y;       // saida

    not(y, a); // porta logica NOT
    
endmodule


