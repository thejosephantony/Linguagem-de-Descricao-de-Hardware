module and2(a, b, y);
    input a, b;     // entradas;
    output y;       // saida

    and(y, a, b);   // porta logica AND
    
endmodule